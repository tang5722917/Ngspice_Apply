INVERSE.CIR - Inverse region operation
* ngspice -a INVERSE.CIR

VCC 2 0 DC 5V ;Supply Voltage 
IB 0 1 DC 1A
Vmess 2 3 dc 0 ;Meassure the E's current
Q1 0 1 3 QC1815   ;2SC1815(Y)

.MODEL QC1815 NPN(IS=1E-14 BF={HFE} xtb=1.7
+                 BR=3.6 VA=100 RB=50 RC=0.76
+                 IK=0.25 CJC=4.8P CJE=18P TF=0.5N TR=20N)
.PARAM HFE = 170

.control
 op
 print ALL > INVERSE_OP.Out
 show Q1  > INVERSE_BJT.Out

 *Output format Control
 DC IB 1uA 1mA 10uA

 set gridstyle=lingrid 
 set xbrushwidth=3   
 set logscale x
 set gnuplot_terminal=png
 gnuplot Inverse I(Vmess) ylimit 0 0.004 xlimit 0 0.001 xlabel 'IB(Q1) A'  ylabel 'IE(Q1) A' title 'Inverse current characteristic' 
 *X轴范围  Y轴范围  X轴名称 Y轴名称  标题名称
.endc
.END