EMF4 - 4 Tr Emitter follower AC sim
* ngspice -a 07_EMF4_AC.CIR

VCC VCC 0 DC +12V
VEE VEE 0 DC -12V
VS 1 0 AC 1V SIN(0 4 1KHZ)
R1 1 2 1K
R2 2 3 47
CF 3 0 10p
R3 6 7 10K
R4 VCC 7 4.7K
R5 9 4 10k
R6 4 VEE 4.7k
R7 10 OUT 47
R8 11 OUT 47
* 自举电容 C1 C2 可使Q1 Q2 的Vcb 交流分量接近0，进而消除米勒效应的影响
C1 7 OUT 33U
C2 8 OUT 33U
RL OUT 0 6K
*<Change> 1 CL OUT 0 <Value>

.INCLUDE ../../../../Spice_Lib/BJT/BJT.mod
.INCLUDE ../../../../Spice_Lib/DIO/DIO.mod

Q1 4 2 5 QA1015
Q2 7 2 8 QC1815
Q3 VCC 6 10 QC2602
Q4 VEE 9 11 QA1114
D1 6 5 DS1588
D2 8 9 DS1588
.control
 run
 op
 *Output format Control
 ac DEC 20 10 100MEG
 let OutDB=DB(VM(OUT)/VM(1))
 wrdata PYTHON_ac1.out.temp ac1.OutDB   ;Print AC data 
.endc
.end