DIODE2.CIR    ;Current Drive
* ngspice -a diode2.cir

Is 0 1 DC 1A 
D1 1 0 DNORM 
.MODEL DNORM D(IS=1E-14)
.PROBE Out = par('V(1)')
.control
 DC Is 1nA 10mA 0.1mA
 *Output format Control
 set gridstyle=lingrid  
 set xbrushwidth=3   
 set gnuplot_terminal=png
 gnuplot DIODE2.CIR Out xlimit 0mA 12mA  ylimit 0.2 0.8V xlabel 'Voltage/V'  ylabel 'Current/A' title 'Current Drive' 
 *X轴范围  Y轴范围  X轴名称 Y轴名称  标题名称
.endc
.END