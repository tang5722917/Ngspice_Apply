CE00.CIR - 1 Transitor circuit
* ngspice -a CE00.CIR
************************
*    Operating  Point
************************
VCC 4 0 DC 12V ;Supply Voltage 
VS 1 0 AC 1 SIN(0 0.01V 1KHZ) ;Inport source
C1 1 2 4.7U
RB 4 2 2MEG
RC 4 3 10K
Q1 3 2 0 QNORM

.MODEL QNORM NPN(IS=1E-14 BF={HFE} xtb=1.7)
.PARAM HFE=100
*.STEP PARAM HFE LIST 50 100 200
.control
 op
 print ALL > CE00_OP.Out
 show Q1  > CE00_BJT.Out

 *Output format Control
 AC DEC 20 10 100K
 let OutDB=DB(VM(3)/VM(1))
 let OutdPH=180/PI*VP(3)
 set gridstyle=lingrid 
 set xbrushwidth=3   
 set logscale x
 set gnuplot_terminal=png
 gnuplot CE00_frequency OutDB ylimit 0 50 xlimit 10 100000 xlabel 'Frequency Hz'  ylabel 'Vo/Vs DB' title 'CE00 frequency characteristic' 
 gnuplot CE00_phase OutdPH ylimit 0 -180 xlimit 10 100000 xlabel 'Frequency Hz'  ylabel 'Phase C' title 'CE00 frequency characteristic' 
 *X轴范围  Y轴范围  X轴名称 Y轴名称  标题名称
.endc
.END