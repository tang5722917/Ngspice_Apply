09_LOWPASS_AC - Butterworth LPF AC  sim
* ngspice -a 09_LOWPASS_AC.CIR

VS 1 0 AC 1

R1 1 2 10K
R2 2 3 10K
C1 2 4 0.02U
C2 3 0 0.01U 
R3 4 OUT 100

RL OUT 0 1MEG
CL OUT 0 300p 

.INCLUDE ../../../Spice_Lib/BJT/BJT.mod
.INCLUDE ../../../Spice_Lib/DIO/DIO.mod

.INCLUDE ../../../Spice_Lib/Module/EMF.mod
X1 3 4 EMF4

.control
 run
 op
 ac DEC 40 10 1Meg
 let OutDB=DB(VM(OUT)/VM(1))
 plot OutDB 
.endc
.END