********** PRE-AMPLIFIER, LOW LEVEL & LOW NOISE   **********
** Product: SS9014
** Package: TO-92
** Terminals: Emitter(1) Base(2) Collector(3)
*BeginSpec
*JV: Ic/Ib=10
*OA: Vce=1
*FB: Vce=1
*VV: Ic/Ib=10
*CB:
*EB:
*ST: Ic/Ib=10
*GB: Vce=10
*EndSpec
*BeginTrace
*JV: 0,1,100.00E-6,.1,1,3,0,0,-1 (27)
*OA: 1,1,100.00E-6,.1,1,3,0,0,-1 (27)
*FB: 0,1,100.00E-6,.1,1,3,0,0,-1 (27)
*VV: 0,1,100.00E-6,.1,1,3,0,0,-1 (27)
*CB: 0,1,.1,50,1,3,0,0,-1 (27)
*EB: 0,1,.1,10,1,3,0,0,-1 (27)
*ST: 0,1,100.00E-6,.1,1,3,0,0,-1 (27)
*GB: 0,1,100.00E-6,.1,1,3,0,0,-1 (27)
*EndTrace
*BeginParam
*IS=10.000E-15 (10.000E-21,1.0000E-6,0)
*BF=100 (1,1.5000E3,0)
*NF=1 (.8,1.2000,0)
*VAF=123 (0,1.0000E3,0)
*IKF=1.1841 (10.000E-3,20,0)
*ISE=4.7863E-15 (0,1,0)
*NE=1.5000 (1,2,0)
*BR=4.7900 (.1,500,0)
*NR=1 (.1,5,0)
*VAR=11.290 (0,1.0000E3,0)
*IKR=.27542 (10.000E-3,20,0)
*ISC=14.454E-15 (0,1,0)
*NC=1.5000 (1,3,0)
*NK=1.1930 (.1,5,0)
*RE=.56 (0,100.00E3,0)
*RB=200 (0,100,0)
*RC=5 (0,100.00E3,0)
*CJE=17.205E-12 (0,1,0)
*VJE=.69059 (.35,1.5000,0)
*MJE=.31934 (.1,1,0)
*CJC=6.2956E-12 (0,1,0)
*VJC=.41642 (.35,1.5000,0)
*MJC=.25595 (.1,1,0)
*FC=.5 (.1,1.5000,0)
*TF=589.46E-12 (0,1,0)
*XTF=10 (0,100.00E3,0)
*VTF=10 (0,100.00E3,0)
*ITF=1 (0,100.00E3,0)
*PTF=0 (0,360,0)
*TR=10.000E-9 (0,1,0)
*EG=1.2415 (.69,5,0)
*XTB=1.8881 (0,100.00E3,0)
*XTI=3 (.1,100.00E3,0)
*EndParam
*DEVICE=SS9014,NPN
* SS9014 NPN model
* created using Model Editor release 10.5.0 on 11/27/08 at 09:05
* The Model Editor is a PSpice product.
.MODEL SS9014 NPN
+ IS=10.000E-15
+ VAF=123             VAR    = 11.29           IKF    = 1.1841             
+ IKF=1.1841             
+ ISE=4.7863E-15         
+ BR=4.7900            NR     = 1               ISE    = 4.7863E-15         
+ VAR=11.290           IKF    = 1.1841             
+ IKR=.27542        NK     = 1.193           RB     = 200                
+ ISC=14.454E-15     NC     = 1.5                
+ NC=1.5000                
+ NK=1.1930           RB     = 200                
+ RE=.56               
+ RB=200                
+ RC=5               CJE    = 1.7205E-11      VJE    = 0.6905907          
+ CJE=17.205E-12      VJE    = 0.6905907          
+ VJE=.69059          
+ MJE=.31934       FC     = 0.5             CJC    = 6.295649E-12       
+ CJC=6.2956E-12       
+ VJC=.41642       MJC    = 0.2559546       TF     = 5.89463E-10        
+ MJC=.25595       TF     = 5.89463E-10        
+ TF=589.46E-12        
+ XTF=10
+ VTF=10
+ ITF=1
+ TR=10.000E-9
+ EG=1.2415          XTI    = 3 
+ XTB=1.8881          EG     = 1.2415          XTI    = 3 
