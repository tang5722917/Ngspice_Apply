06_EMF3_THD - EMF3 - 3 Tr emitter follower
* ngspice -a 02_EMF3_THD.CIR

VCC 6 0 DC 5V ;Supply Voltage 
VEE 10 0 DC -5V
VSS 1 0 AC 1 SIN(0 {VIN} 1KHZ)
*Vs 1 0 AC 1V sin(0 {VIN} 20KHz)

R1 1 2 47
R2 6 5 100
R3 4 10 1K
R4 4 9 100
R5 6 7 39
R6 8 out 75
RL out 0 6k
CL out 0 20p 
D1 5 3 DS1588
Q1 3 2 4 QC1815 
Q2 10 9 8 QA1114
Q3 8 3 7 QA1114

*<Change> 1 RL 8 out 6k  ;RL = 6k

*<Change> 2 RL 8 0 75  ;RL = 75

.INCLUDE ../../../Spice_Lib/BJT/BJT.mod
.INCLUDE ../../../Spice_Lib/DIO/DIO.mod
.PARAM VIN = 1

.tran 5us 1ms 0 5u 
.probe I(Q1,c) I(Q3,e)
.control
 alterparam VIN = 1
 run
 let Out_Q1x2.5 = Q1:c#branch * 2.5 
 plot Out_Q1x2.5 Q3:e#branch
.endc
.END