STAGE2A_with_boost.CIR - Common emitter+common collector
* ngspice -a STAGE2A_with_boost.CIR

VCC 10 0 DC 12V ;Supply Voltage 
Vs 1 0 AC 1V sin(0 {VIN} 1KHz)
*Vs 1 0 AC 1V sin(0 {VIN} 20KHz)
R0 1 0 22k
C1 1 2 10U
R1 2 3 2.2K
R2 3 6 4.7K
R3 9 10 10K
R4 9 4 10K
C2 9 5 47U      ;with boost capacitor
R5 5 6 910
R6 6 0 100
R7 5 7 470
C3 7 8 220U
RL 8 0 6K
Q1 4 3 0 QC2240
Q2 10 4 5 QC1815

.INCLUDE ../../../Spice_Lib/BJT/BJT.mod
.PARAM VIN = 1

*.TRAN 10US 1MS

.control
 run
 op
 print ALL > STAGE2A_OP.Out
 show Q1 Q2 > STAGE2A_BJT.Out
 *Output format Control
 ac DEC 20 10 10MEG
 let OutDB=DB(VM(8)/VM(1))
 write STAGE2A-sweepAC1.out OutDB
 wrdata STAGE2A_ac2.out ac1.OutDB
.endc
.END