DIODE1.CIR    ;Current Drive
* ngspice -a diode2.cir

Is 0 1 DC 1A 
D1 1 0 DNORM 
.DC Is 1nA 10mA 0.1mA
.MODEL DNORM D(IS=1E-14)
.PROBE 

.control
 
 run 
 set gridstyle=lingrid  ;坐标轴
 set xbrushwidth=3   ;线宽
 plot v(1) ylimit 0 2V xlimit 0mA 1mA  xlabel Current_Drive ylabel Voltage title 1.2  
 *X轴范围  Y轴范围  X轴名称 Y轴名称  标题名称
.endc
.END