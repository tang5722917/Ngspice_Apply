STAGE2_THD.CIR - Common emitter+common collector
* stage2b - NPN + PNP
* ngspice -a STAGE2B_AC_CF.CIR

VCC 11 0 DC 12V ;Supply Voltage 
Vs 2 0 AC 1V sin(0 {VIN} 1KHz)

R1 1 0 100K
R2 1 2 470
C1 2 3 3.3U
C2 3 0 56p
R3 11 3 100K
R4 3 0 120K
R5 3 4 100
Q1 5 4 6 QC2240  ;2SC2240
Q2 7 5 11 QA1015 ;2SA1015

CF 5 7 5P

R6 11 5 4.7K
R7 6 7 220
R8 7 0 1K
R9 7 8 220
C3 8 9 220U
RL 9 0 6K

.INCLUDE ../../../Spice_Lib/BJT/BJT.mod
.PARAM VIN = 0.1

.control
 *Output format Control
 ac DEC 20 10 100MEG
 let OutDB=DB(VM(9)/VM(2))
 wrdata STAGE2A_ac1.out ac1.OutDB
 plot ac1.OutDB
.endc
.END