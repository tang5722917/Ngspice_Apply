04_STAGE2B_AC_CF - Common emitter+common collector
* stage2b - NPN + PNP
* ngspice -a 04_STAGE2B_AC_CF.CIR

VCC 11 0 DC 12V ;Supply Voltage 
Vs 1 0 AC 1V sin(0 {VIN} 1KHz)

R1 1 0 100K
R2 1 2 470
C1 2 3 3.3U
C2 3 0 56p
R3 11 3 100K
R4 3 0 120K
R5 3 4 100
Q1 5_Q 4 6 QC2240  ;2SC2240
Q2 7 5 11 QA1015 ;2SA1015
*CF 5 7 22P 
*<Change> 1 CF 5 7 <Value> ;Difference value of CF

R6 11 5 4.7K

R7 6 7 220
R8 7 0 1K
R9 7 8 220
C3 8 9 220U
RL 9 0 6K

V_Q1_Ic 5 5_Q DC 0
.PARAM VIN = 1
.INCLUDE ../../../../Spice_Lib/BJT/BJT.mod

.control
 run
 op
 *Output format Control
 ac DEC 20 10 100MEG
 let OutDB=DB(VM(9)/VM(2))
 wrdata PYTHON_ac1.out.temp ac1.OutDB   ;Print AC data 
*plot OutDB
.endc
.END
