01_TRANSFORMER ST7 - 01_TRANSFORMER ST71
* ngspice -a 01_TRANSFORMER_ST71.CIR
V1 100 0 ac 1
Rs 100 1 50
X1 1 0 2 0 3 ST71 
*<Change> 1 RL 2 3 <Value>

.SUBCKT ST71 1 2 3 4 5
R1 1 6 51
C1 1 2 400p 
L1 6 2 1.2
L2 7 4 0.3
L3 4 8 0.3
C2 3 5 400p 
K12 L1 L2 0.9992
K13 L1 L3 0.9992
K23 L2 L3 0.9995
R2 7 3 27.5
R3 8 5 27.5
.ENDS 
.control
 run
 op
 *Output format Control
 ac DEC 50 10 200k
 let OutDB=DB(VM(3)/VM(1))
 wrdata PYTHON_ac1.out.temp ac1.OutDB   ;Print AC data 
.endc
.END
