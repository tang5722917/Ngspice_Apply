01_SQUARE_WAVE - Square wave Oscillator 
* ngspice -a 01_SQUARE_WAVE.CIR

VCC VCC 0 DC 12V  ;Supply Voltage 
VEE VEE 0 DC -12V

R1 NI 0 10k
R2 OUT NI 47K
R3 OUT INV 47k
C1 INV 0 0.01U IC=1V
X1 NI INV OUT CMP VCC VEE OPAMP3

.SUBCKT OPAMP3 NI INV OUT CMP VCC VEE
R1 VCC 1 30K
R2 CMP VEE 3.9K
R3 VCC OUT 2.2K
Q1 CMP NI 1 QA872A
Q2 VEE INV 1 QA872A
Q3 OUT CMP VEE QC1815 
.ENDS


.INCLUDE ../../../Spice_Lib/BJT/BJT.mod
.OP
.tran 2us 1ms 0 2U UIC 

.control
run
plot V(OUT) V(NI) V(INV)
.endc
.END