CE00A.CIR - 1 Transitor circuit
* ngspice -a CE01.CIR
************************
*    BIAS TYPE no.
*    ARAM HFE = 120 170 240
************************

VCC 5 0 DC 5V ;Supply Voltage 
VS 1 0 AC 1V SIN(0 0.05V 1KHZ) ;Import source
C1 1 2 3.3U
RB1 2 3 4.7K
RB2 4 3 220K
Q1 4 3 0 QC1815   ;2SC1815(Y)
RC 5 4 1.5K
R1 4 6 220
C2 6 7 1.5U
RL1 7 0 1MEG
CL 7 0 300P

*C3 6 8 220U
*RL2 8 0 6K
*.FOUR 1KHz V(8)

.MODEL QC1815 NPN(IS=1E-14 BF={HFE} xtb=1.7
+                 BR=3.6 VA=100 RB=50 RC=0.76
+                 IK=0.25 CJC=4.8P CJE=18P TF=0.5N TR=20N)
.PARAM HFE = 50
.tran 10us 2ms 0 10us 

.control
 *.STEP PARAM HFE LIST 120 170 240
 altermod QC1815 BF = 120
 run
 write HFE-sweep.out V(6)
 set appendwrite
 altermod QC1815 BF = 170
 run
 write HFE-sweep.out V(6)
 set appendwrite
 altermod QC1815 BF = 240
 run
 write HFE-sweep.out V(6)
 set appendwrite

 *Output format Control
 set gridstyle=lingrid
 set xbrushwidth=3   
 set gnuplot_terminal=png
 wrdata outfile.out tran1.V(6) tran2.V(6) tran3.V(6)
 *gnuplot CE01_HFE_120 tran1.V(6) tran2.V(6) tran3.V(6) ;ylimit 1 4 xlimit 0 0.002 xlabel 'Frequency Hz'  ylabel 'Vo/Vs DB' title 'CE00 frequency characteristic' 
 *X轴范围  Y轴范围  X轴名称 Y轴名称  标题名称
.endc
.END