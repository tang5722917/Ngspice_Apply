CASCODE - Wide freq range amp
* ngspice -a  CASCODE.CIR

VCC VCC 0 DC +12V
VEE VEE 0 DC -12V
VS 1 0 AC 1V PWL ( 0 0.0 1N 0.8
+ 0.5U 0.8 0.501U -0.8 1U -0.8
+          1.001U 0.8 1.2U 0.8)
R1 1 2 200
R2 4 5 97
R3 6 5 97
R4 5 VEE 3.9K 
R5 7 0 200 
R6 VCC 3 300
R7 VCC 8 300

.INCLUDE ../../../Spice_Lib/BJT/BJT.mod
.INCLUDE ../../../Spice_Lib/DIO/DIO.mod
Q1 3  2  4  2SC1775
Q2 8  7  6  2SC1775
Q3 9  11 8  QA1015
Q4 10 11 3  QA1015
Q5 17 9  16 QC1815
C1 10  17  0.01U 
D1 9   15  DS1588 
R8 15 VEE  150 
R9 16 VEE  150
R10 11 12  47
D2 VCC 14   DS1588
D3 14  13   DS1588  
D4 13  12   DS1588
D5 10  19   DS1588
D6 19  18   DS1588
D7 18  17   DS1588
Q6 VCC 10 20  QC1815
Q7 VEE 17 22  QA1015
R11 12 VEE 10K 
R12 20 21  33 
R13 21 22  33
R14 21 2   2K
R15 21 OUT  51
CL  OUT 0   20P   


.control
run
op
tran 0.01U 1.2U 0 0.01U
 *Output format Control
*ac DEC 20 10 100MEG
*let OutDB=DB(VM(OUT)/VM(1))
*plot OutDB
plot V(OUT) V(1)
 *wrdata PYTHON_ac1.out.temp ac1.OutDB   ;Print AC data 
.endc
.end
